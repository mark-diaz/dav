module miniALU (
    input [3:0] op1,
    input [3:0] op2, 
    input operation,
    input sign,
    output [19:0] result
    );

    always_comb begin
        

    end
endmodule